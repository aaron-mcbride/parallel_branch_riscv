`ifndef __STACK_SV__
`define __STACK_SV__

// Stack module
module stack #(
  parameter int size = 32,
  parameter type data_type = logic [31:0]
) (
  input logic clk,
  input logic rst,
  input logic 
)

`endif // __STACK_SV__
`include "common.sv"

`ifndef __HZD_UNIT_SV__
`define __HZD_UNIT_SV__

module hzd_unit (
  input logic clk,
  input bool rst,
  input bool en,

);

`endif // __HZD_UNIT_SV__